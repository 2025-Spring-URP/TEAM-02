// Copyright (c) 2024 Sungkyunkwan University
// All rights reserved
// Author: YongSeong Lim <xidid430rr@gmail.com>
// Description:

module SAL_FIFO
#(



)
(





);

//AXI_Interface
//FIFO






endmodule