// 1 ) Decoder - TLP / DLLP check
// 2 ) 

// NAK_Scheduled