// Timer
// Next_RCV_SEQ
// NAK_SCHEDULED