module CRC_CHECKER
#(

)
(

);



endmodule