module _DLL_DLCMSM(
	input wire clk,
	



);

endmodule