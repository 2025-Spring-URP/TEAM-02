// Timer
// NAK_SCHEDULED


module _DLL_DLLP_Generator
#(

)
(
    // -------------------------------------------------------
    //                    DLCMSM
    // -------------------------------------------------------
    input   wire     [1:0]                          DLCM_state,         // LINK_UP, LINK_DOWN

);

endmodule