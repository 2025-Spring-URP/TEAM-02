// 

module _DLL_Arbitor
#(

)
(
    // -------------------------------------------------------
    //                    DLCMSM
    // -------------------------------------------------------
    input   wire                                    DL_up,







);

endmodule