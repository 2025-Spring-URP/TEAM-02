// SEQ + LCRC 붙이기.
