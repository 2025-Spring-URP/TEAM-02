// Receive_TLP_FIFO!

module DLL_TOP (

    output  wire                             dll2tl_data_en_o;
);


endmodule
